`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2022/10/14 10:04:15
// Design Name: 
// Module Name: CP0
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

// д�ؽ׶�
 module CP0(
	input			reset,
	input           clock,
    
    input           Overflow,
    input           Divide_zero,
    input           Reserved_instruction,
    input           Mfc0,           // ��Ȩָ��
    input           Mtc0,
    input           Break,
    input           Syscall,
    input           Eret,
    input [5:0]     ExternalInterrupt,
    input           backFromEret,//��һ��ָ����Eret

    input [31:0]    PC,
    input [4:0]     rd,
    input [31:0]    rt_value,     //д������ 
    output reg      cp0_wen,
    output reg[31:0] cp0_data_out,
    output reg[31:0] cp0_pc_out
    );
    wire [4:0] causeExcCode;
    reg wen;
    reg [31:0] cp0[0:31];   // cp0����32���Ĵ���
    reg status_IE;          // �ж�����
    reg [1:0] status_KSU;   // 
    
    //�ⲿ�ж��������ڲ��ж�
    assign causeExcCode = (ExternalInterrupt[0]===1'b1) ? 5'b00000 :   // �����ⲿ�ж�
                          (ExternalInterrupt[1]===1'b1) ? 5'b01101 :   // button S1
                          (ExternalInterrupt[2]===1'b1) ? 5'b01110 :   // button S2
                          (ExternalInterrupt[3]===1'b1) ? 5'b01111 :   // button S3
                          (ExternalInterrupt[4]===1'b1) ? 5'b10000 :   // button S4
                          (ExternalInterrupt[5]===1'b1) ? 5'b10001 :   // button S5
                          (Syscall===1'b1) ? 5'b01000 :                // ϵͳ���� syscall
                          (Divide_zero===1'b1) ? 5'b00111:             // �������
                          (Break===1'b1) ? 5'b01001 :                  // ���Զϵ�ָ�� break
                          (Reserved_instruction===1'b1) ? 5'b01010 :   // ����ָ��,cpuִ�е�һ��δ�����ָ��
                          (Overflow===1'b1) ?  5'b01100 :              // ����������з�������Ӽ����
                          5'b11111;  
    integer i;                
    always @(negedge clock) begin
        if(reset) begin
            for(i=0;i<32;i=i+1)
                cp0[i] = 0; 
            cp0[12][0] = 1'b1;
            cp0[12][15:10] = 6'b111111;
        end
        wen = (causeExcCode!=5'b11111)&&(!backFromEret)&&cp0[12][0];//cp0[12][0]���ж���Ч
        cp0_wen = wen||Eret;  
        if(Mtc0===1'b1) begin
            cp0[rd] = rt_value;
        end else if(Eret===1'b1) begin
            // Step1. �ָ� CP0.Status.KSU ��ԭʼֵ
            cp0[12][4:3] = status_KSU;
            // Step2. �ָ� CP0.Status.IE
            //cp0[12][0] = status_IE;
            cp0[12][0] = 1'b1;
            // Step3. PC<-EPC
            cp0_pc_out = cp0[14];
        end else if(wen===1'b1) begin // �ж���Ӧ�Ĺ���
            // Step1. ���� CP0.Status.IE
            // status_IE = cp0[12][0];
            // Step2. CP0.Status.IE<-0 �������жϣ�
            cp0[12][0] = 1'b0;
            // Step3. ���� CP0.Status.KSU
            status_KSU = cp0[12][4:3];
            // Step4. CP0.Status.KSU<-0�������Ĳ㣩,KSU-CPU ��Ȩ����0 Ϊ���ļ���2 Ϊ�û���
            cp0[12][4:3] = 2'b00;
            // Step5. �����жϡ��쳣�źŻ�ִ�е��� Break �� SysCall ָ���д CP0.Cause.ExcCode
            cp0[13][6:2] = causeExcCode;
            // Step6. EPC<-PC�����淵�ص�ַ��
            cp0[14] = PC;
            // Step7. PC<-�жϴ��������ڵ�ַ�������жϺ��쳣ֻ��һ����ڵ�ַ��32'h0x0000F500��
            cp0_pc_out = 32'h0000F500;
        end
    end 
    
    always @(*) begin
        if(reset) begin // ��ʼ����cp0�Ĵ���ȫ����ֵ0
            cp0_data_out = 32'h00000000;
        end else begin
            if(Mfc0===1'b1) begin
                cp0_data_out = cp0[rd];
            end 
        end
    end
    
endmodule
